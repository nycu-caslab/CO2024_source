/*
*  Description
*    - alu has two input operand a and b.
*    - alu executes different operation over input a and b based on input s
*    - alu outputs final result to y
*/

module alu(
    input signed [3:0] a,
    input signed [3:0] b,
    input [2:0] s,
    output reg signed [3:0] y
); 
    
    // TODO: implement your 4bits ALU design here and using your own fulladder module in this module
    // For testbench verifying, do not modify input and output pin
    
endmodule

